library verilog;
use verilog.vl_types.all;
entity Task3_16071005_vlg_vec_tst is
end Task3_16071005_vlg_vec_tst;
