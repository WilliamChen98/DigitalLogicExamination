library verilog;
use verilog.vl_types.all;
entity TenthProject_vlg_sample_tst is
    port(
        clk             : in     vl_logic;
        clr             : in     vl_logic;
        rst             : in     vl_logic;
        sel             : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end TenthProject_vlg_sample_tst;
