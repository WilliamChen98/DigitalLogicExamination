module divider(ind,outkd,outmd);
	input[3:0]ind;
	output reg[3:0]outkd,outmd;
	always @ (ind)
		case(ind)
			4'd0:outkd = ind;
			4'd1:outkd = ind;
			4'd2:outkd = ind;
			4'd3:outkd = ind;
			4'd4:outkd = ind;
			4'd5:outkd = ind;
			4'd6:outkd = ind;
			4'd7:outkd = ind;
			4'd8:outkd = ind;
			4'd9:outkd = ind;
			4'd10:outmd = ind;
			4'd11:outmd = ind;
			4'd12:outmd = ind;
			4'd13:outmd = ind;
			4'd14:outmd = ind;
			4'd15:outmd = ind;
			default:begin outkd = outkd;outmd = outmd; end
		endcase
endmodule