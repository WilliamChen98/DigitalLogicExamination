library verilog;
use verilog.vl_types.all;
entity Task3_16071005_vlg_check_tst is
    port(
        count           : in     vl_logic_vector(2 downto 0);
        sampler_rx      : in     vl_logic
    );
end Task3_16071005_vlg_check_tst;
