library verilog;
use verilog.vl_types.all;
entity count_dis_vlg_vec_tst is
end count_dis_vlg_vec_tst;
