library verilog;
use verilog.vl_types.all;
entity Counter_2421_16071005 is
    port(
        clk             : in     vl_logic;
        Q               : out    vl_logic_vector(3 downto 0);
        z               : out    vl_logic
    );
end Counter_2421_16071005;
