library verilog;
use verilog.vl_types.all;
entity xl_reciver_vlg_vec_tst is
end xl_reciver_vlg_vec_tst;
