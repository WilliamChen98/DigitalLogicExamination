library verilog;
use verilog.vl_types.all;
entity xl_generate_vlg_vec_tst is
end xl_generate_vlg_vec_tst;
