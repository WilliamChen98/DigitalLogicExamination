library verilog;
use verilog.vl_types.all;
entity scaner_vlg_vec_tst is
end scaner_vlg_vec_tst;
