library verilog;
use verilog.vl_types.all;
entity FifthProject_vlg_vec_tst is
end FifthProject_vlg_vec_tst;
