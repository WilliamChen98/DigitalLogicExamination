library verilog;
use verilog.vl_types.all;
entity Second_vlg_vec_tst is
end Second_vlg_vec_tst;
