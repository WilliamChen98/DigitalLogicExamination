library verilog;
use verilog.vl_types.all;
entity NinthProject_00_vlg_vec_tst is
end NinthProject_00_vlg_vec_tst;
