library verilog;
use verilog.vl_types.all;
entity Demux8Way_vlg_vec_tst is
end Demux8Way_vlg_vec_tst;
