library verilog;
use verilog.vl_types.all;
entity Register_8_vlg_vec_tst is
end Register_8_vlg_vec_tst;
