library verilog;
use verilog.vl_types.all;
entity TenthProject_vlg_vec_tst is
end TenthProject_vlg_vec_tst;
