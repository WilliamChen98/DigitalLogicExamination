library verilog;
use verilog.vl_types.all;
entity check_vlg_vec_tst is
end check_vlg_vec_tst;
