library verilog;
use verilog.vl_types.all;
entity xl_generate_vlg_check_tst is
    port(
        dout            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end xl_generate_vlg_check_tst;
