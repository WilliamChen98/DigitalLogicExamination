library verilog;
use verilog.vl_types.all;
entity Fifth_vlg_vec_tst is
end Fifth_vlg_vec_tst;
