library verilog;
use verilog.vl_types.all;
entity price_count_vlg_vec_tst is
end price_count_vlg_vec_tst;
