library verilog;
use verilog.vl_types.all;
entity testoften_vlg_vec_tst is
end testoften_vlg_vec_tst;
