library verilog;
use verilog.vl_types.all;
entity Counter_2421_16071005_vlg_vec_tst is
end Counter_2421_16071005_vlg_vec_tst;
