library verilog;
use verilog.vl_types.all;
entity Tenth_vlg_vec_tst is
end Tenth_vlg_vec_tst;
