library verilog;
use verilog.vl_types.all;
entity Eleventhproject_vlg_vec_tst is
end Eleventhproject_vlg_vec_tst;
