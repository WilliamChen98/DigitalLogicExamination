library verilog;
use verilog.vl_types.all;
entity Eleventh_vlg_vec_tst is
end Eleventh_vlg_vec_tst;
