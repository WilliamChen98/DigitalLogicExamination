library verilog;
use verilog.vl_types.all;
entity Counter_2421_16071005_vlg_check_tst is
    port(
        Q               : in     vl_logic_vector(3 downto 0);
        z               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Counter_2421_16071005_vlg_check_tst;
